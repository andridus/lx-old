module token

pub struct Token {
	pub mut:
	 typ string
	 literal string
}