module docs

pub const (
	local_function_desc = 'The local functions should be defined in the context of the module before they\ncan be used anywhere in the module.'
	local_function_url = 'https://github.com/andridus/lx/wiki/Refer%C3%AAncia-da-Linguagem#funcoes-locais'

)