module parser

import compiler_v.types
import compiler_v.ast

pub fn (p Parser) node_string_left(node string) ast.NodeLeft {
	return ast.NodeLeft(node)
}

pub fn (p Parser) node_left(node ast.Node) ast.NodeLeft {
	return ast.NodeLeft(node)
}

pub fn (p Parser) node(meta ast.Meta, left ast.NodeLeft, nodes []ast.Node) ast.Node {
	kind := match left {
		string {
			match left {
				'defmodule' {
					ast.NodeKind(ast.Module{})
				}
				'def' {
					ast.NodeKind(ast.Ast{
						lit: 'def'
					})
				}
				'__aliases__' {
					ast.NodeKind(ast.Alias{})
				}
				'.' {
					ast.NodeKind(ast.Ast{
						lit: '.'
					})
				}
				'__block__' {
					ast.NodeKind(ast.Ast{
						lit: 'block'
					})
				}
				else {
					ast.NodeKind(ast.Nil{})
				}
			}
		}
		ast.Node {
			left.kind
		}
	}
	return ast.Node{
		left: left
		kind: kind
		meta: meta
		nodes: nodes
	}
}

pub fn (p Parser) node_function(meta ast.Meta, left ast.NodeLeft, nodes []ast.Node, ty ast.Function) ast.Node {
	return ast.Node{
		left: left
		kind: ast.NodeKind(ty)
		meta: meta
		nodes: nodes
	}
}

pub fn (p Parser) node_function_caller(meta ast.Meta, left ast.NodeLeft, nodes []ast.Node, ty ast.FunctionCaller) ast.Node {
	return ast.Node{
		left: left
		kind: ast.NodeKind(ty)
		meta: meta
		nodes: nodes
	}
}

pub fn (p Parser) node_var(meta ast.Meta, left string, nodes []ast.Node) ast.Node {
	return ast.Node{
		left: ast.NodeLeft(left)
		kind: ast.NodeKind(ast.Ast{
			lit: 'var'
		})
		meta: meta
		nodes: nodes
	}
}

pub fn (p Parser) node_assign(meta ast.Meta, ident string, node ast.Node) ast.Node {
	return ast.Node{
		left: ast.NodeLeft('=')
		kind: ast.NodeKind(ast.Ast{
			lit: 'assign'
		})
		meta: meta
		nodes: [p.node_var(meta, ident, []), node]
	}
}

pub fn (p Parser) node_atom(mut meta ast.Meta, atom string) ast.Node {
	meta.put_ti(types.atom_ti)
	return ast.Node{
		left: ast.NodeLeft(atom)
		kind: ast.NodeKind(ast.Atom{})
		meta: meta
	}
}

pub fn (p Parser) node_string(mut meta ast.Meta, str string) ast.Node {
	meta.put_ti(types.string_ti)
	return ast.Node{
		left: ast.NodeLeft(str)
		kind: ast.NodeKind(ast.String{})
		meta: meta
	}
}

pub fn (p Parser) node_integer(mut meta ast.Meta, val int) ast.Node {
	meta.put_ti(types.integer_ti)
	return ast.Node{
		left: ast.NodeLeft(val.str())
		kind: ast.NodeKind(ast.Integer{})
		meta: meta
	}
}

pub fn (p Parser) node_float(mut meta ast.Meta, val f64) ast.Node {
	meta.put_ti(types.float_ti)
	return ast.Node{
		left: ast.NodeLeft(val.str())
		kind: ast.NodeKind(ast.Float{})
		meta: meta
	}
}

pub fn (p Parser) node_tuple(meta ast.Meta, nodes []ast.Node) ast.Node {
	return ast.Node{
		kind: ast.NodeKind(ast.Tuple{})
		meta: meta
		nodes: nodes
	}
}

pub fn (p Parser) node_list(meta ast.Meta, nodes []ast.Node) ast.Node {
	return ast.Node{
		kind: ast.NodeKind(ast.List{})
		meta: meta
		nodes: nodes
	}
}

pub fn (p Parser) node_atomic(atom string) ast.Node {
	return ast.Node{
		left: ast.NodeLeft(atom)
		kind: ast.NodeKind(ast.Atomic{})
		nodes: []
	}
}

pub fn (p Parser) node_default() ast.Node {
	return ast.Node{
		left: ast.NodeLeft('default')
		kind: ast.NodeKind(ast.Atomic{})
		nodes: []
	}
}

pub fn (p Parser) meta() ast.Meta {
	return ast.Meta{
		line: p.tok.line_nr
		inside_parens: p.inside_parens
	}
}
